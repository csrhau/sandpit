library ieee;
use ieee.std_logic_1164.all;

package three_multiple_types is
  type three_state is (SAccept, S1, S2); 
end package three_multiple_types;
