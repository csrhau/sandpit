library ieee;
use ieee.std_logic_1164.all;

entity test_slv is 
end test_slv;

architecture behavioural of test_slv is

begin
  process
  begin

    wait;
  end process;
end behavioural;
